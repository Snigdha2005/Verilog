module tb_mux4;
reg d0;
reg d1;
reg d2;
reg d3;
reg sel1;
reg sel2;
wire Data_out;
mux4 namexyz1(d0,d1,d2,d3,sel1,sel2,Data_out);
initial
begin
	$dumpfile("mux4_out.vcd");
	$dumpvars(0,tb_mux4);
	d0=0;
	d1=0;
	d2=0;
	d3=0;
	sel1=0;
	sel2=0;
	#10;

	d0=0;	d1=0;	d2=0;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=0;	d2=0;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=0;	d2=0;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=0;	d1=0;	d2=0;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=0;	d1=0;	d2=0;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=0;	d2=0;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=0;	d2=0;	d3=1;	sel1=1;	sel2=1;	#10;
	d0=0;	d1=0;	d2=1;	d3=0;	sel1=0;	sel2=0;	#10;
	d0=0;	d1=0;	d2=1;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=0;	d2=1;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=0;	d2=1;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=0;	d1=0;	d2=1;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=0;	d1=0;	d2=1;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=0;	d2=1;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=0;	d2=1;	d3=1;	sel1=1;	sel2=1;	#10;
	d0=0;	d1=1;	d2=0;	d3=0;	sel1=0;	sel2=0;	#10;
	d0=0;	d1=1;	d2=0;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=1;	d2=0;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=1;	d2=0;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=0;	d1=1;	d2=0;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=0;	d1=1;	d2=0;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=1;	d2=0;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=1;	d2=0;	d3=1;	sel1=1;	sel2=1;	#10;
	d0=0;	d1=1;	d2=1;	d3=0;	sel1=0;	sel2=0;	#10;
	d0=0;	d1=1;	d2=1;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=1;	d2=1;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=1;	d2=1;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=0;	d1=1;	d2=1;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=0;	d1=1;	d2=1;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=0;	d1=1;	d2=1;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=0;	d1=1;	d2=1;	d3=1;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=0;	d2=0;	d3=0;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=0;	d2=0;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=0;	d2=0;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=0;	d2=0;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=0;	d2=0;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=0;	d2=0;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=0;	d2=0;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=0;	d2=0;	d3=1;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=0;	d2=1;	d3=0;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=0;	d2=1;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=0;	d2=1;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=0;	d2=1;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=0;	d2=1;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=0;	d2=1;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=0;	d2=1;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=0;	d2=1;	d3=1;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=1;	d2=0;	d3=0;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=1;	d2=0;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=1;	d2=0;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=1;	d2=0;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=1;	d2=0;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=1;	d2=0;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=1;	d2=0;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=1;	d2=0;	d3=1;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=1;	d2=1;	d3=0;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=1;	d2=1;	d3=0;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=1;	d2=1;	d3=0;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=1;	d2=1;	d3=0;	sel1=1;	sel2=1;	#10;
	d0=1;	d1=1;	d2=1;	d3=1;	sel1=0;	sel2=0;	#10;
	d0=1;	d1=1;	d2=1;	d3=1;	sel1=0;	sel2=1;	#10;
	d0=1;	d1=1;	d2=1;	d3=1;	sel1=1;	sel2=0;	#10;
	d0=1;	d1=1;	d2=1;	d3=1;	sel1=1;	sel2=1;	#10;
end
endmodule
